*** SPICE deck for cell logic_CONTROL_II{sch} from library SIPO_register
*** Created on Sun Dec 10, 2023 18:42:14
*** Last revised on Thu Dec 28, 2023 20:57:05
*** Written on Thu Dec 28, 2023 20:57:12 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include /home/miqueasgamero/my_files/VLSI/Models/models.txt

*** SUBCIRCUIT SIPO_register__ffsr_sOK FROM CELL ffsr_sOK{sch}
.SUBCKT SIPO_register__ffsr_sOK CLK Q Qn R S
** GLOBAL gnd
** GLOBAL vdd
Mnmos-4@0 Qn Q gnd nmos-4@0_b NMOS L=0.6U W=1.8U
Mnmos-4@1 Qn S net@6 nmos-4@1_b NMOS L=0.6U W=1.8U
Mnmos-4@2 net@6 CLK gnd nmos-4@2_b NMOS L=0.6U W=1.8U
Mnmos-4@3 Q Qn gnd nmos-4@3_b NMOS L=0.6U W=1.8U
Mnmos-4@4 Q R net@31 nmos-4@4_b NMOS L=0.6U W=1.8U
Mnmos-4@5 net@31 CLK gnd nmos-4@5_b NMOS L=0.6U W=1.8U
Mpmos-4@0 vdd S net@11 pmos-4@0_b PMOS L=0.6U W=3U
Mpmos-4@1 vdd CLK net@11 pmos-4@1_b PMOS L=0.6U W=3U
Mpmos-4@2 net@11 Q Qn pmos-4@2_b PMOS L=0.6U W=3U
Mpmos-4@6 vdd R net@21 pmos-4@6_b PMOS L=0.6U W=3U
Mpmos-4@7 vdd CLK net@21 pmos-4@7_b PMOS L=0.6U W=3U
Mpmos-4@8 net@21 Qn Q pmos-4@8_b PMOS L=0.6U W=3U
.ENDS SIPO_register__ffsr_sOK

*** SUBCIRCUIT SIPO_register__inv FROM CELL inv{sch}
.SUBCKT SIPO_register__inv in out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out in gnd gnd NMOS L=0.6U W=1.8U
Mpmos@0 vdd in out vdd PMOS L=0.6U W=3U
.ENDS SIPO_register__inv

*** SUBCIRCUIT SIPO_register__nand FROM CELL nand{sch}
.SUBCKT SIPO_register__nand A B out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out A net@10 gnd NMOS L=0.6U W=1.8U
Mnmos@1 net@10 B gnd gnd NMOS L=0.6U W=1.8U
Mpmos@0 vdd A out vdd PMOS L=0.6U W=3U
Mpmos@1 vdd B out vdd PMOS L=0.6U W=3U
.ENDS SIPO_register__nand

*** SUBCIRCUIT SIPO_register__and FROM CELL and{sch}
.SUBCKT SIPO_register__and A B out
** GLOBAL gnd
** GLOBAL vdd
Xinv@0 net@0 out SIPO_register__inv
Xnand@0 A B net@0 SIPO_register__nand
.ENDS SIPO_register__and

*** SUBCIRCUIT SIPO_register__logic_OUTPUTs FROM CELL logic_OUTPUTs{sch}
.SUBCKT SIPO_register__logic_OUTPUTs ACK CK Q0 Q0_ Q1 Q1_ TG
** GLOBAL gnd
** GLOBAL vdd
Xand@0 Q1 Q0_ ACK SIPO_register__and
Xand@1 Q0 Q1_ CK SIPO_register__and
Xand@2 Q0 Q1 TG SIPO_register__and
.ENDS SIPO_register__logic_OUTPUTs

*** SUBCIRCUIT SIPO_register__and3 FROM CELL and3{sch}
.SUBCKT SIPO_register__and3 A B C out
** GLOBAL gnd
** GLOBAL vdd
Mnmos-4@0 net@1 A net@9 nmos-4@0_b NMOS L=0.6U W=1.8U
Mnmos-4@1 net@9 B net@10 nmos-4@1_b NMOS L=0.6U W=1.8U
Mnmos-4@2 net@10 C gnd nmos-4@2_b NMOS L=0.6U W=1.8U
Mnmos-4@4 out net@1 gnd nmos-4@4_b NMOS L=0.6U W=1.8U
Mpmos-4@0 vdd A net@1 pmos-4@0_b PMOS L=0.6U W=3U
Mpmos-4@1 vdd B net@1 pmos-4@1_b PMOS L=0.6U W=3U
Mpmos-4@2 vdd C net@1 pmos-4@2_b PMOS L=0.6U W=3U
Mpmos-4@4 vdd net@1 out pmos-4@4_b PMOS L=0.6U W=3U
.ENDS SIPO_register__and3

*** SUBCIRCUIT SIPO_register__nor FROM CELL nor{sch}
.SUBCKT SIPO_register__nor A B out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out A gnd gnd NMOS L=0.6U W=1.8U
Mnmos@1 out B gnd gnd NMOS L=0.6U W=1.8U
Mpmos@0 vdd A net@20 vdd PMOS L=0.6U W=3U
Mpmos@1 net@20 B out vdd PMOS L=0.6U W=3U
.ENDS SIPO_register__nor

*** SUBCIRCUIT SIPO_register__or FROM CELL or{sch}
.SUBCKT SIPO_register__or A B out
** GLOBAL gnd
** GLOBAL vdd
Xinv@0 net@0 out SIPO_register__inv
Xnor@0 A B net@0 SIPO_register__nor
.ENDS SIPO_register__or

*** SUBCIRCUIT SIPO_register__logic_R1 FROM CELL logic_R1{sch}
.SUBCKT SIPO_register__logic_R1 EN Q0 Q0_ Q1 R1
** GLOBAL gnd
** GLOBAL vdd
Xand3@0 EN Q0_ Q1 net@16 SIPO_register__and3
Xand@0 net@1 Q0 net@14 SIPO_register__and
Xinv@0 EN net@1 SIPO_register__inv
Xor@0 net@14 net@16 R1 SIPO_register__or
.ENDS SIPO_register__logic_R1

*** SUBCIRCUIT SIPO_register__logic_S0R0 FROM CELL logic_S0R0{sch}
.SUBCKT SIPO_register__logic_S0R0 EN Q1 R0 S0 SYN
** GLOBAL gnd
** GLOBAL vdd
Xand@12 EN net@114 net@129 SIPO_register__and
Xand@13 EN Q1 net@127 SIPO_register__and
Xinv@2 SYN net@114 SIPO_register__inv
Xinv@3 EN R0 SIPO_register__inv
Xor@3 net@127 net@129 S0 SIPO_register__or
.ENDS SIPO_register__logic_S0R0

*** SUBCIRCUIT SIPO_register__and4 FROM CELL and4{sch}
.SUBCKT SIPO_register__and4 A B C D out
** GLOBAL gnd
** GLOBAL vdd
Mnmos-4@0 net@1 A net@9 nmos-4@0_b NMOS L=0.6U W=1.8U
Mnmos-4@1 net@9 B net@10 nmos-4@1_b NMOS L=0.6U W=1.8U
Mnmos-4@2 net@10 C net@11 nmos-4@2_b NMOS L=0.6U W=1.8U
Mnmos-4@3 net@11 D gnd nmos-4@3_b NMOS L=0.6U W=1.8U
Mnmos-4@4 out net@1 gnd nmos-4@4_b NMOS L=0.6U W=1.8U
Mpmos-4@0 vdd A net@1 pmos-4@0_b PMOS L=0.6U W=3U
Mpmos-4@1 vdd B net@1 pmos-4@1_b PMOS L=0.6U W=3U
Mpmos-4@2 vdd C net@1 pmos-4@2_b PMOS L=0.6U W=3U
Mpmos-4@3 vdd D net@1 pmos-4@3_b PMOS L=0.6U W=3U
Mpmos-4@4 vdd net@1 out pmos-4@4_b PMOS L=0.6U W=3U
.ENDS SIPO_register__and4

*** SUBCIRCUIT SIPO_register__logic_S1 FROM CELL logic_S1{sch}
.SUBCKT SIPO_register__logic_S1 EN Q0_ Q1_ S1 SYN
** GLOBAL gnd
** GLOBAL vdd
Xand3@1 SYN net@43 Q0_ net@0 SIPO_register__and3
Xand4@0 net@75 EN Q0_ Q1_ net@61 SIPO_register__and4
Xinv@0 SYN net@75 SIPO_register__inv
Xinv@1 EN net@43 SIPO_register__inv
Xor@0 net@61 net@0 S1 SIPO_register__or
.ENDS SIPO_register__logic_S1

.global gnd vdd

*** TOP LEVEL CELL: logic_CONTROL_II{sch}
VPulse@0 CLK gnd DC=1V pulse 0 5V 0ns 200ps 200ps 5ns 10ns
VPulse@1 SYN gnd DC=1V pulse 0 5V 20ns 200ps 200ps 10ns 100ns
VPulse@2 EN gnd DC=1V pulse 0 5V 50ns 200ps 200ps 20ns 100ns
Xffsr_s@0 CLK Q0 net@28 net@12 net@15 SIPO_register__ffsr_sOK
Xffsr_s@1 CLK Q1 net@22 net@9 net@6 SIPO_register__ffsr_sOK
Xlogic_OU@0 ACK CK Q0 net@28 Q1 net@22 TG SIPO_register__logic_OUTPUTs
Xlogic_R1@0 EN Q0 net@28 Q1 net@9 SIPO_register__logic_R1
Xlogic_S0@0 EN Q1 net@12 net@15 SYN SIPO_register__logic_S0R0
Xlogic_S1@0 EN net@28 net@22 net@6 SYN SIPO_register__logic_S1

* Spice Code nodes in cell cell 'logic_CONTROL_II{sch}'
vdd vdd 0 DC 5 
.tran 100n
.END
